
module decode_jump_inst(
    input logic [31:0] instruction_code,
    output logic [4:0] rd,
    output logic [4:0] rs1,
    output logic [20:0] imm,
    output logic [1:0] jump_control
);



endmodule
